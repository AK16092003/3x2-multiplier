module multiply(x,y,q);

	input [2:0] x; 
	input [1:0] y;
	output [4:0] Q;

	assign Q[0] = (x[0] && y[0]);
	assign Q[1] = ((x[1]&&y[0])^(x[0]&&y[1]));
	assign Q[2] = ((x[1] && y[0] && x[0] && y[1])^(x[2]&&y[0]))^(x[1]&&y[1]);
    assign Q[3] = (x[2]&&y[1])^((x[1]&&y[0]&& x[0] && y[1])&&((x[2]&&y[0])||(x[1]&&y[1]))|| (x[2]&&y[0]&&x[1]&&y[1]));
	assign Q[4] = (x[2]&&y[1]) && ((x[1]&&y[0]&& x[0] && y[1])&&((x[2]&&y[0])||(x[1]&&y[1]))|| (x[2]&&y[0]&&x[1]&&y[1]));
	
endmodule